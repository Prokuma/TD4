module ROM (
	input [3:0] ADDR,
	output reg [7:0] COMMAND
);

always @* begin
	case (ADDR)
		4'b0000: COMMAND <= 8'b10110111;
		4'b0001: COMMAND <= 8'b00000001;
		4'b0010: COMMAND <= 8'b11100001;
		4'b0011: COMMAND <= 8'b00000001;
		4'b0100: COMMAND <= 8'b11100011;
		4'b0101: COMMAND <= 8'b10110110;
		4'b0110: COMMAND <= 8'b00000001;
		4'b0111: COMMAND <= 8'b11100110;
		4'b1000: COMMAND <= 8'b00000001;
		4'b1001: COMMAND <= 8'b11101000;
		4'b1010: COMMAND <= 8'b10110000;
		4'b1011: COMMAND <= 8'b10110100;
		4'b1100: COMMAND <= 8'b00000001;
		4'b1101: COMMAND <= 8'b11101010;
		4'b1110: COMMAND <= 8'b10111000;
		4'b1111: COMMAND <= 8'b11111111;
	endcase
end

endmodule