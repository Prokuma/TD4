module TD4(
	input CLK,
	input [3:0] IN,
	output [3:0] OUT
);

wire [1:0] SEL;
wire [3:0] LOAD, REGA_OUT, REGB_OUT, ADDR, SEL_OUT, IM, ALU_OUT;
wire [7:0] COMMAND;
reg CFLAG_IN;
wire CFLAG_OUT;

REG REG_A(.CLK(CLK), .LOAD(LOAD[0]), .IN(ALU_OUT), .CNT(0), .OUT(REGA_OUT));
REG REG_B(.CLK(CLK), .LOAD(LOAD[1]), .IN(ALU_OUT), .CNT(0), .OUT(REGB_OUT));
REG REG_O(.CLK(CLK), .LOAD(LOAD[2]), .IN(ALU_OUT), .CNT(0), .OUT(OUT));
REG REG_P(.CLK(CLK), .LOAD(LOAD[3]), .IN(ALU_OUT), .CNT(1), .OUT(ADDR));

SELECTOR SELECTOR (.REGA(REGA_OUT), .REGB(REGB_OUT), .IN(IN), .SEL(SEL), .OUT(SEL_OUT));

ROM ROM(.ADDR(ADDR), .COMMAND(COMMAND));

ALU ALU(.INPUT(SEL_OUT), .IM(IM), .OUTPUT(ALU_OUT), .CFLAG(CFLAG_OUT));

DECODER DECODER(.COMMAND(COMMAND), .CFLAG(CFLAG_IN), .IM(IM), .LOAD(LOAD), .SEL(SEL));

always @(posedge CLK) begin
	CFLAG_IN <= CFLAG_OUT;
end

endmodule